module fault_detector (
    input   NS_RED,
    input   NS_YELLOW,
    input   NS_GREEN,

    input   EW_RED,
    input   EW_YELLOW,
    input   EW_GREEN
    
);

endmodule