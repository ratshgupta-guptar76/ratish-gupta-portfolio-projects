module traffic_controller (
    input clk,
    output dbg,
);

    
endmodule